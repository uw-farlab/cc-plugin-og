netcdf bad_variable {
dimensions:
	N_MEASUREMENTS = 66 ;
	N_BINS = 20 ;
	traj_strlen = 22 ;
variables:
	double time(N_MEASUREMENTS) ;
		time:_FillValue = -9999.9 ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:comment = "Measured or calculated time at each point in the time-series" ;
		time:long_name = "Time" ;
		time:observation_type = "measured" ;
		time:ioos_category = "Time" ;
		time:coordinates = "lat_uv lon_uv time_uv" ;
		time:units = "seconds since 1990-01-01T00:00:00+00:00" ;
		time:calendar = "gregorian" ;
	double depth(N_MEASUREMENTS, N_BINS) ;
		depth:_FillValue = NaN ;
		depth:axis = "Z" ;
		depth:accuracy = "n/a" ;
		depth:long_name = "Depth" ;
		depth:observation_type = "calculated" ;
		depth:platform = "platform" ;
		depth:precision = "n/a" ;
		depth:resolution = "n/a" ;
		depth:positive = "down" ;
		depth:reference_datum = "sea-surface" ;
		depth:standard_name = "depth" ;
		depth:units = "m" ;
		depth:valid_max = 2000. ;
		depth:valid_min = 0. ;
		depth:ioos_category = "Location" ;
		depth:colorBarMaximum = 2000. ;
		depth:colorBarMinimum = 0. ;
		depth:colorBarPalette = "OceanDepth" ;
		depth:instrument = "instrument_altimeter" ;
		depth:comment = "Native glider sensor name" ;
		depth:coordinates = "lat_uv lon_uv time_uv" ;
	double echogram_sv(N_MEASUREMENTS, N_BINS) ;
		echogram_sv:_FillValue = NaN ;
		echogram_sv:units = "1" ;
		echogram_sv:long_name = "Volume backscattering strength" ;
		echogram_sv:colorBarMinimum = -80. ;
		echogram_sv:colorBarMaximum = -30. ;
		echogram_sv:colorBarPalette = "EK80" ;
		echogram_sv:comment = "dimensionless units (dB re 1 m-1)" ;
		echogram_sv:ioos_category = "Other" ;
		echogram_sv:standard_name = "acoustic_volume_backscattering_strength_in_sea_water" ;
		echogram_sv:platform = "platform" ;
		echogram_sv:observation_type = "measured" ;
		echogram_sv:coordinates = "lat_uv lon_uv time_uv" ;
	double lat(N_MEASUREMENTS) ;
		lat:_FillValue = NaN ;
		lat:axis = "Y" ;
		lat:comment = "Interpolated latitude at each point in the time-series" ;
		lat:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lat:long_name = "Precise Latitude" ;
		lat:observation_type = "measured" ;
		lat:platform = "platform" ;
		lat:reference = "WGS84" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_max = 90. ;
		lat:valid_min = -90. ;
		lat:ioos_category = "Location" ;
		lat:colorBarMaximum = 90. ;
		lat:colorBarMinimum = -90. ;
		lat:coordinates = "lat_uv lon_uv time_uv" ;
	double lon(N_MEASUREMENTS) ;
		lon:_FillValue = NaN ;
		lon:axis = "X" ;
		lon:comment = "Interpolated longitude at each point in the time-series." ;
		lon:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lon:long_name = "Precise Longitude" ;
		lon:observation_type = "measured" ;
		lon:platform = "platform" ;
		lon:reference = "WGS84" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_max = 180. ;
		lon:valid_min = -180. ;
		lon:ioos_category = "Location" ;
		lon:colorBarMaximum = 180. ;
		lon:colorBarMinimum = -180. ;
		lon:coordinates = "lat_uv lon_uv time_uv" ;
	double lat_uv ;
		lat_uv:_FillValue = -9999.9 ;
		lat_uv:long_name = "Depth-Averaged Latitude" ;
		lat_uv:valid_max = 90. ;
		lat_uv:observation_type = "calculated" ;
		lat_uv:colorBarMaximum = 90. ;
		lat_uv:ioos_category = "Location" ;
		lat_uv:standard_name = "latitude" ;
		lat_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		lat_uv:units = "degrees_north" ;
		lat_uv:platform = "platform" ;
		lat_uv:valid_min = -90. ;
		lat_uv:colorBarMinimum = -90. ;
	double lon_uv ;
		lon_uv:_FillValue = -9999.9 ;
		lon_uv:long_name = "Depth-Averaged Longitude" ;
		lon_uv:valid_max = 180. ;
		lon_uv:observation_type = "calculated" ;
		lon_uv:colorBarMaximum = 180. ;
		lon_uv:ioos_category = "Location" ;
		lon_uv:standard_name = "longitude" ;
		lon_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		lon_uv:units = "degrees_east" ;
		lon_uv:platform = "platform" ;
		lon_uv:valid_min = -180. ;
		lon_uv:colorBarMinimum = -180. ;
	double time_uv ;
		time_uv:_FillValue = -9999.9 ;
		time_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		time_uv:long_name = "Depth-Averaged Time" ;
		time_uv:observation_type = "calculated" ;
		time_uv:standard_name = "time" ;
		time_uv:ioos_category = "Time" ;
		time_uv:units = "seconds since 1990-01-01T00:00:00+00:00" ;
		time_uv:calendar = "gregorian" ;
	int profile_id ;
		profile_id:_FillValue = -999 ;
		profile_id:comment = "Sequential profile number within the trajectory.  This value is unique in each file that is part of a single trajectory/deployment." ;
		profile_id:long_name = "Profile ID" ;
		profile_id:valid_max = 2147483647 ;
		profile_id:valid_min = 0 ;
		profile_id:cf_role = "profile_id" ;
		profile_id:ioos_category = "Identifier" ;
		profile_id:coordinates = "lat_uv lon_uv time_uv" ;
	double profile_lat ;
		profile_lat:_FillValue = -9999.9 ;
		profile_lat:long_name = "Profile Latitude" ;
		profile_lat:valid_max = 90. ;
		profile_lat:observation_type = "calculated" ;
		profile_lat:colorBarMaximum = 90. ;
		profile_lat:ioos_category = "Location" ;
		profile_lat:standard_name = "latitude" ;
		profile_lat:comment = "Value is interpolated to provide an estimate of the latitude at the mid-point of the profile" ;
		profile_lat:units = "degrees_north" ;
		profile_lat:platform = "platform" ;
		profile_lat:valid_min = -90. ;
		profile_lat:colorBarMinimum = -90. ;
		profile_lat:coordinates = "lat_uv lon_uv time_uv" ;
	double profile_lon ;
		profile_lon:_FillValue = -9999.9 ;
		profile_lon:long_name = "Profile Longitude" ;
		profile_lon:valid_max = 180. ;
		profile_lon:observation_type = "calculated" ;
		profile_lon:colorBarMaximum = 180. ;
		profile_lon:ioos_category = "Location" ;
		profile_lon:standard_name = "longitude" ;
		profile_lon:comment = "Value is interpolated to provide an estimate of the longitude at the mid-point of the profile" ;
		profile_lon:units = "degrees_east" ;
		profile_lon:platform = "platform" ;
		profile_lon:valid_min = -180. ;
		profile_lon:colorBarMinimum = -180. ;
		profile_lon:coordinates = "lat_uv lon_uv time_uv" ;
	double profile_time ;
		profile_time:_FillValue = -9999.9 ;
		profile_time:long_name = "Profile Time" ;
		profile_time:observation_type = "calculated" ;
		profile_time:ioos_category = "Time" ;
		profile_time:standard_name = "time" ;
		profile_time:comment = "Timestamp corresponding to the mid-point of the profile" ;
		profile_time:platform = "platform" ;
		profile_time:coordinates = "lat_uv lon_uv time_uv" ;
		profile_time:units = "seconds since 1990-01-01T00:00:00+00:00" ;
		profile_time:calendar = "gregorian" ;
	double u ;
		u:_FillValue = -9999.9 ;
		u:long_name = "Depth-Averaged Eastward Sea Water Velocity" ;
		u:valid_max = 10. ;
		u:observation_type = "calculated" ;
		u:colorBarMaximum = 0.5 ;
		u:ioos_category = "Currents" ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		u:units = "m.s-1" ;
		u:platform = "platform" ;
		u:valid_min = -10. ;
		u:colorBarMinimum = -0.5 ;
		u:coordinates = "lon_uv lat_uv time_uv" ;
	double v ;
		v:_FillValue = -9999.9 ;
		v:long_name = "Depth-Averaged Northward Sea Water Velocity" ;
		v:valid_max = 10. ;
		v:observation_type = "calculated" ;
		v:colorBarMaximum = 0.5 ;
		v:ioos_category = "Currents" ;
		v:standard_name = "northward_sea_water_velocity" ;
		v:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		v:units = "m.s-1" ;
		v:platform = "platform" ;
		v:valid_min = -10. ;
		v:colorBarMinimum = -0.5 ;
		v:coordinates = "lon_uv lat_uv time_uv" ;
	int platform ;
		platform:_FillValue = -999 ;
		platform:type = "platform" ;
		platform:long_name = "G507 Slocum Glider" ;
		platform:ioos_category = "Identifier" ;
		platform:wmo_id = 4802989 ;
		platform:comment = "Teledyne Webb Research Slocum G2 Glider" ;
		platform:id = 4802989 ;
		platform:instrument = "instrument_ctd,instrument_acoustics" ;
		platform:coordinates = "lat_uv lon_uv time_uv" ;
	int instrument_ctd ;
		instrument_ctd:_FillValue = 0 ;
		instrument_ctd:calibration_report = "n/a" ;
		instrument_ctd:long_name = "Seabird WEBB pumped glider conductivity, temperature, depth sensor" ;
		instrument_ctd:factory_calibrated = "y" ;
		instrument_ctd:type = "instrument" ;
		instrument_ctd:serial_number = "712-9221" ;
		instrument_ctd:comment = "Slocum Glider UAF G507 -- pumped CTD" ;
		instrument_ctd:user_calibrated = "n/a" ;
		instrument_ctd:platform = "platform" ;
		instrument_ctd:make_model = "Seabird Slocum Glider Payload CTD" ;
		instrument_ctd:calibration_date = "2017" ;
		instrument_ctd:coordinates = "lat_uv lon_uv time_uv" ;
	char trajectory(traj_strlen) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:long_name = "Trajectory/Deployment Name" ;
		trajectory:comment = "A trajectory is a single deployment of a glider and may span multiple data files." ;
		trajectory:ioos_category = "Identifier" ;
		trajectory:coordinates = "lat_uv lon_uv time_uv" ;

// global attributes:
		:Conventions = "OG-1.0,CF-1.10" ;
		:date_created = "2024-03-22T01:21:12Z" ;
		:featureType = "trajectoryProfile" ;
		:cdm_data_type = "trajectory" ;
		:comment = "UAF G507 Glider deployment in the North Pacific Ocean (March 2024)" ;
		:format_version = "IOOS_Glider_NetCDF_v2.0.nc" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:keywords = "Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:license = "This data may be redistributed and used without restriction." ;
		:Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:metadata_link = "https://gliders.ioos.us/erddap/info/unit_507-20240304T0000/index.html" ;
		:platform_type = "Slocum Glider" ;
		:processing_level = "Dataset taken from glider native file format and is provided as is with no expressed or implied assurance of quality assurance or quality control." ;
		:project = "AOOS Gliders in Support of Fisheries Management" ;
		:references = "https://www.uaf.edu/cfos/" ;
		:source = "Observational data from a profiling glider" ;
		:standard_name_vocabulary = "Standard Name Table (v84a)" ;
		:summary = "UAF G507 Glider deployment in the North Pacific Ocean (March 2024)" ;
		:title = "G507 Slocum Glider Dataset (March 2024)" ;
		:acknowledgement = "This work was supported by funding from NOAA/IOOS/AOOS." ;
		:contributor_email = "sldanielson@alaska.edu" ;
		:contributor_name = "Seth Danielson" ;
		:contributor_role = "Principal Investigator" ;
		:contributor_url = "https://www.uaf.edu/cfos/people/faculty/detail/seth-danielson.php" ;
		:creator_email = "hank.stats@alaska.edu" ;
		:creator_name = "Hank Statscewich" ;
		:creator_url = "https://uaf.edu/cfos/people/research-staff-and-post-docs/detail/hank-statscewich.php" ;
		:institution = "The University of Alaska Fairbanks College of Fisheries and Ocean Sciences" ;
		:ioos_regional_association = "aoos" ;
		:naming_authority = "edu.alaska" ;
		:platform_tags = "portal:25,axds:portal:25:tag:Gliders,axds:dashboard:glider:EcoMetrics Dashboard" ;
		:publisher_email = "dmac@aoos.org" ;
		:publisher_name = "AOOS Glider Observatory" ;
		:publisher_url = "https://aoos.org" ;
		:sea_name = "North Pacific Ocean" ;
		:support_email = "dmac@aoos.org,ioos.glider.data@noaa.gov,ioos.glider.data@noaa.gov" ;
		:support_name = "aoos,ioos,noaa" ;
		:support_role = "fiscal,fiscal,fiscal" ;
		:support_type = "ra,federal,federal" ;
		:wmo_id = 4802989 ;
		:geospatial_lat_min = 59.83922 ;
		:geospatial_lat_max = 59.8421 ;
		:geospatial_lon_min = -149.47692 ;
		:geospatial_lon_max = -149.47529 ;
		:geospatial_bounds = "POLYGON ((59.842100 -149.476920, 59.842100 -149.475290, 59.839220 -149.475290, 59.839220 -149.476920, 59.842100 -149.476920))" ;
		:geospatial_vertical_min = 1.407026 ;
		:geospatial_vertical_max = 200.89151 ;
		:geospatial_vertical_units = "m" ;
		:time_coverage_start = "2024-03-13T20:46:09Z" ;
		:time_coverage_end = "2024-03-13T21:07:11Z" ;
		:time_coverage_duration = "P0DT0H21M2.478820864S" ;
		:date_issued = "2024-03-22T01:21:12Z" ;
		:date_modified = "2024-03-22T01:21:12Z" ;
		:history = "2024-03-22T01:21:12Z - Created with the GUTILS package: https://github.com/SECOORA/GUTILS" ;
		:id = "unit_507-20240304T0000" ;
data:

 time = 1079210769.3107, 1079210823.87811, 1079210843.11444, 
    1079210861.31677, 1079210880.47821, 1079210899.73987, 1079210917.97824, 
    1079210937.21442, 1079210955.51129, 1079210974.69778, 1079210993.93704, 
    1079211012.13187, 1079211031.35004, 1079211050.59244, 1079211068.82413, 
    1079211088.08414, 1079211107.33133, 1079211125.5705, 1079211144.8013, 
    1079211163.98578, 1079211182.2316, 1079211201.48706, 1079211219.71576, 
    1079211238.93393, 1079211258.19183, 1079211276.35315, 1079211295.48285, 
    1079211314.59253, 1079211333.70746, 1079211351.82446, 1079211370.90518, 
    1079211389.98102, 1079211409.22284, 1079211427.41132, 1079211446.62744, 
    1079211465.88534, 1079211484.12485, 1079211503.35443, 1079211521.64407, 
    1079211540.86838, 1079211560.11118, 1079211578.29343, 1079211597.53802, 
    1079211616.76047, 1079211635.00482, 1079211654.228, 1079211673.47107, 
    1079211691.68076, 1079211710.84463, 1079211730.09985, 1079211748.30179, 
    1079211767.5639, 1079211785.86224, 1079211805.05545, 1079211824.28693, 
    1079211842.45563, 1079211861.7066, 1079211880.91977, 1079211899.16354, 
    1079211918.40506, 1079211937.64313, 1079211955.86728, 1079211975.10645, 
    1079211994.28238, 1079212012.52759, 1079212031.78952 ;

 depth =
  143.891510009766, 146.891510009766, 149.891510009766, 152.891510009766, 
    155.891510009766, 158.891510009766, 161.891510009766, 164.891510009766, 
    167.891510009766, 170.891510009766, 173.891510009766, 176.891510009766, 
    179.891510009766, 182.891510009766, 185.891510009766, 188.891510009766, 
    191.891510009766, 194.891510009766, 197.891510009766, 200.891510009766,
  138.106964111328, 141.106964111328, 144.106964111328, 147.106964111328, 
    150.106964111328, 153.106964111328, 156.106964111328, 159.106964111328, 
    162.106964111328, 165.106964111328, 168.106964111328, 171.106964111328, 
    174.106964111328, 177.106964111328, 180.106964111328, 183.106964111328, 
    186.106964111328, 189.106964111328, 192.106964111328, 195.106964111328,
  134.5859375, 137.5859375, 140.5859375, 143.5859375, 146.5859375, 
    149.5859375, 152.5859375, 155.5859375, 158.5859375, 161.5859375, 
    164.5859375, 167.5859375, 170.5859375, 173.5859375, 176.5859375, 
    179.5859375, 182.5859375, 185.5859375, 188.5859375, 191.5859375,
  130.897232055664, 133.897232055664, 136.897232055664, 139.897232055664, 
    142.897232055664, 145.897232055664, 148.897232055664, 151.897232055664, 
    154.897232055664, 157.897232055664, 160.897232055664, 163.897232055664, 
    166.897232055664, 169.897232055664, 172.897232055664, 175.897232055664, 
    178.897232055664, 181.897232055664, 184.897232055664, 187.897232055664,
  127.3203125, 130.3203125, 133.3203125, 136.3203125, 139.3203125, 
    142.3203125, 145.3203125, 148.3203125, 151.3203125, 154.3203125, 
    157.3203125, 160.3203125, 163.3203125, 166.3203125, 169.3203125, 
    172.3203125, 175.3203125, 178.3203125, 181.3203125, 184.3203125,
  123.771347045898, 126.771347045898, 129.771347045898, 132.771347045898, 
    135.771347045898, 138.771347045898, 141.771347045898, 144.771347045898, 
    147.771347045898, 150.771347045898, 153.771347045898, 156.771347045898, 
    159.771347045898, 162.771347045898, 165.771347045898, 168.771347045898, 
    171.771347045898, 174.771347045898, 177.771347045898, 180.771347045898,
  120.25032043457, 123.25032043457, 126.25032043457, 129.25032043457, 
    132.25032043457, 135.25032043457, 138.25032043457, 141.25032043457, 
    144.25032043457, 147.25032043457, 150.25032043457, 153.25032043457, 
    156.25032043457, 159.25032043457, 162.25032043457, 165.25032043457, 
    168.25032043457, 171.25032043457, 174.25032043457, 177.25032043457,
  116.393951416016, 119.393951416016, 122.393951416016, 125.393951416016, 
    128.393951416016, 131.393951416016, 134.393951416016, 137.393951416016, 
    140.393951416016, 143.393951416016, 146.393951416016, 149.393951416016, 
    152.393951416016, 155.393951416016, 158.393951416016, 161.393951416016, 
    164.393951416016, 167.393951416016, 170.393951416016, 173.393951416016,
  116.393951416016, 119.393951416016, 122.393951416016, 125.393951416016, 
    128.393951416016, 131.393951416016, 134.393951416016, 137.393951416016, 
    140.393951416016, 143.393951416016, 146.393951416016, 149.393951416016, 
    152.393951416016, 155.393951416016, 158.393951416016, 161.393951416016, 
    164.393951416016, 167.393951416016, 170.393951416016, 173.393951416016,
  112.956756591797, 115.956756591797, 118.956756591797, 121.956756591797, 
    124.956756591797, 127.956756591797, 130.956756591797, 133.956756591797, 
    136.956756591797, 139.956756591797, 142.956756591797, 145.956756591797, 
    148.956756591797, 151.956756591797, 154.956756591797, 157.956756591797, 
    160.956756591797, 163.956756591797, 166.956756591797, 169.956756591797,
  109.407775878906, 112.407775878906, 115.407775878906, 118.407775878906, 
    121.407775878906, 124.407775878906, 127.407775878906, 130.407775878906, 
    133.407775878906, 136.407775878906, 139.407775878906, 142.407775878906, 
    145.407775878906, 148.407775878906, 151.407775878906, 154.407775878906, 
    157.407775878906, 160.407775878906, 163.407775878906, 166.407775878906,
  105.830856323242, 108.830856323242, 111.830856323242, 114.830856323242, 
    117.830856323242, 120.830856323242, 123.830856323242, 126.830856323242, 
    129.830856323242, 132.830856323242, 135.830856323242, 138.830856323242, 
    141.830856323242, 144.830856323242, 147.830856323242, 150.830856323242, 
    153.830856323242, 156.830856323242, 159.830856323242, 162.830856323242,
  102.36572265625, 105.36572265625, 108.36572265625, 111.36572265625, 
    114.36572265625, 117.36572265625, 120.36572265625, 123.36572265625, 
    126.36572265625, 129.36572265625, 132.36572265625, 135.36572265625, 
    138.36572265625, 141.36572265625, 144.36572265625, 147.36572265625, 
    150.36572265625, 153.36572265625, 156.36572265625, 159.36572265625,
  98.9564666748047, 101.956466674805, 104.956466674805, 107.956466674805, 
    110.956466674805, 113.956466674805, 116.956466674805, 119.956466674805, 
    122.956466674805, 125.956466674805, 128.956466674805, 131.956466674805, 
    134.956466674805, 137.956466674805, 140.956466674805, 143.956466674805, 
    146.956466674805, 149.956466674805, 152.956466674805, 155.956466674805,
  95.2677764892578, 98.2677764892578, 101.267776489258, 104.267776489258, 
    107.267776489258, 110.267776489258, 113.267776489258, 116.267776489258, 
    119.267776489258, 122.267776489258, 125.267776489258, 128.267776489258, 
    131.267776489258, 134.267776489258, 137.267776489258, 140.267776489258, 
    143.267776489258, 146.267776489258, 149.267776489258, 152.267776489258,
  91.7746887207031, 94.7746887207031, 97.7746887207031, 100.774688720703, 
    103.774688720703, 106.774688720703, 109.774688720703, 112.774688720703, 
    115.774688720703, 118.774688720703, 121.774688720703, 124.774688720703, 
    127.774688720703, 130.774688720703, 133.774688720703, 136.774688720703, 
    139.774688720703, 142.774688720703, 145.774688720703, 148.774688720703,
  88.3933868408203, 91.3933868408203, 94.3933868408203, 97.3933868408203, 
    100.39338684082, 103.39338684082, 106.39338684082, 109.39338684082, 
    112.39338684082, 115.39338684082, 118.39338684082, 121.39338684082, 
    124.39338684082, 127.39338684082, 130.39338684082, 133.39338684082, 
    136.39338684082, 139.39338684082, 142.39338684082, 145.39338684082,
  84.9282379150391, 87.9282379150391, 90.9282379150391, 93.9282379150391, 
    96.9282379150391, 99.9282379150391, 102.928237915039, 105.928237915039, 
    108.928237915039, 111.928237915039, 114.928237915039, 117.928237915039, 
    120.928237915039, 123.928237915039, 126.928237915039, 129.928237915039, 
    132.928237915039, 135.928237915039, 138.928237915039, 141.928237915039,
  84.9282379150391, 87.9282379150391, 90.9282379150391, 93.9282379150391, 
    96.9282379150391, 99.9282379150391, 102.928237915039, 105.928237915039, 
    108.928237915039, 111.928237915039, 114.928237915039, 117.928237915039, 
    120.928237915039, 123.928237915039, 126.928237915039, 129.928237915039, 
    132.928237915039, 135.928237915039, 138.928237915039, 141.928237915039,
  81.2395477294922, 84.2395477294922, 87.2395477294922, 90.2395477294922, 
    93.2395477294922, 96.2395477294922, 99.2395477294922, 102.239547729492, 
    105.239547729492, 108.239547729492, 111.239547729492, 114.239547729492, 
    117.239547729492, 120.239547729492, 123.239547729492, 126.239547729492, 
    129.239547729492, 132.239547729492, 135.239547729492, 138.239547729492,
  77.718505859375, 80.718505859375, 83.718505859375, 86.718505859375, 
    89.718505859375, 92.718505859375, 95.718505859375, 98.718505859375, 
    101.718505859375, 104.718505859375, 107.718505859375, 110.718505859375, 
    113.718505859375, 116.718505859375, 119.718505859375, 122.718505859375, 
    125.718505859375, 128.718505859375, 131.718505859375, 134.718505859375,
  74.4210357666016, 77.4210357666016, 80.4210357666016, 83.4210357666016, 
    86.4210357666016, 89.4210357666016, 92.4210357666016, 95.4210357666016, 
    98.4210357666016, 101.421035766602, 104.421035766602, 107.421035766602, 
    110.421035766602, 113.421035766602, 116.421035766602, 119.421035766602, 
    122.421035766602, 125.421035766602, 128.421035766602, 131.421035766602,
  71.2632904052734, 74.2632904052734, 77.2632904052734, 80.2632904052734, 
    83.2632904052734, 86.2632904052734, 89.2632904052734, 92.2632904052734, 
    95.2632904052734, 98.2632904052734, 101.263290405273, 104.263290405273, 
    107.263290405273, 110.263290405273, 113.263290405273, 116.263290405273, 
    119.263290405273, 122.263290405273, 125.263290405273, 128.263290405273,
  68.1055374145508, 71.1055374145508, 74.1055374145508, 77.1055374145508, 
    80.1055374145508, 83.1055374145508, 86.1055374145508, 89.1055374145508, 
    92.1055374145508, 95.1055374145508, 98.1055374145508, 101.105537414551, 
    104.105537414551, 107.105537414551, 110.105537414551, 113.105537414551, 
    116.105537414551, 119.105537414551, 122.105537414551, 125.105537414551,
  64.7521820068359, 67.7521820068359, 70.7521820068359, 73.7521820068359, 
    76.7521820068359, 79.7521820068359, 82.7521820068359, 85.7521820068359, 
    88.7521820068359, 91.7521820068359, 94.7521820068359, 97.7521820068359, 
    100.752182006836, 103.752182006836, 106.752182006836, 109.752182006836, 
    112.752182006836, 115.752182006836, 118.752182006836, 121.752182006836,
  61.5664825439453, 64.5664825439453, 67.5664825439453, 70.5664825439453, 
    73.5664825439453, 76.5664825439453, 79.5664825439453, 82.5664825439453, 
    85.5664825439453, 88.5664825439453, 91.5664825439453, 94.5664825439453, 
    97.5664825439453, 100.566482543945, 103.566482543945, 106.566482543945, 
    109.566482543945, 112.566482543945, 115.566482543945, 118.566482543945,
  58.4087371826172, 61.4087371826172, 64.4087371826172, 67.4087371826172, 
    70.4087371826172, 73.4087371826172, 76.4087371826172, 79.4087371826172, 
    82.4087371826172, 85.4087371826172, 88.4087371826172, 91.4087371826172, 
    94.4087371826172, 97.4087371826172, 100.408737182617, 103.408737182617, 
    106.408737182617, 109.408737182617, 112.408737182617, 115.408737182617,
  58.4087371826172, 61.4087371826172, 64.4087371826172, 67.4087371826172, 
    70.4087371826172, 73.4087371826172, 76.4087371826172, 79.4087371826172, 
    82.4087371826172, 85.4087371826172, 88.4087371826172, 91.4087371826172, 
    94.4087371826172, 97.4087371826172, 100.408737182617, 103.408737182617, 
    106.408737182617, 109.408737182617, 112.408737182617, 115.408737182617,
  55.2789306640625, 58.2789306640625, 61.2789306640625, 64.2789306640625, 
    67.2789306640625, 70.2789306640625, 73.2789306640625, 76.2789306640625, 
    79.2789306640625, 82.2789306640625, 85.2789306640625, 88.2789306640625, 
    91.2789306640625, 94.2789306640625, 97.2789306640625, 100.278930664062, 
    103.278930664062, 106.278930664062, 109.278930664062, 112.278930664062,
  52.1491317749023, 55.1491317749023, 58.1491317749023, 61.1491317749023, 
    64.1491317749023, 67.1491317749023, 70.1491317749023, 73.1491317749023, 
    76.1491317749023, 79.1491317749023, 82.1491317749023, 85.1491317749023, 
    88.1491317749023, 91.1491317749023, 94.1491317749023, 97.1491317749023, 
    100.149131774902, 103.149131774902, 106.149131774902, 109.149131774902,
  49.2708282470703, 52.2708282470703, 55.2708282470703, 58.2708282470703, 
    61.2708282470703, 64.2708282470703, 67.2708282470703, 70.2708282470703, 
    73.2708282470703, 76.2708282470703, 79.2708282470703, 82.2708282470703, 
    85.2708282470703, 88.2708282470703, 91.2708282470703, 94.2708282470703, 
    97.2708282470703, 100.27082824707, 103.27082824707, 106.27082824707,
  46.0571899414062, 49.0571899414062, 52.0571899414062, 55.0571899414062, 
    58.0571899414062, 61.0571899414062, 64.0571899414062, 67.0571899414062, 
    70.0571899414062, 73.0571899414062, 76.0571899414062, 79.0571899414062, 
    82.0571899414062, 85.0571899414062, 88.0571899414062, 91.0571899414062, 
    94.0571899414062, 97.0571899414062, 100.057189941406, 103.057189941406,
  43.0950546264648, 46.0950546264648, 49.0950546264648, 52.0950546264648, 
    55.0950546264648, 58.0950546264648, 61.0950546264648, 64.0950546264648, 
    67.0950546264648, 70.0950546264648, 73.0950546264648, 76.0950546264648, 
    79.0950546264648, 82.0950546264648, 85.0950546264648, 88.0950546264648, 
    91.0950546264648, 94.0950546264648, 97.0950546264648, 100.095054626465,
  39.7975769042969, 42.7975769042969, 45.7975769042969, 48.7975769042969, 
    51.7975769042969, 54.7975769042969, 57.7975769042969, 60.7975769042969, 
    63.7975769042969, 66.7975769042969, 69.7975769042969, 72.7975769042969, 
    75.7975769042969, 78.7975769042969, 81.7975769042969, 84.7975769042969, 
    87.7975769042969, 90.7975769042969, 93.7975769042969, 96.7975769042969,
  36.6677780151367, 39.6677780151367, 42.6677780151367, 45.6677780151367, 
    48.6677780151367, 51.6677780151367, 54.6677780151367, 57.6677780151367, 
    60.6677780151367, 63.6677780151367, 66.6677780151367, 69.6677780151367, 
    72.6677780151367, 75.6677780151367, 78.6677780151367, 81.6677780151367, 
    84.6677780151367, 87.6677780151367, 90.6677780151367, 93.6677780151367,
  33.56591796875, 36.56591796875, 39.56591796875, 42.56591796875, 
    45.56591796875, 48.56591796875, 51.56591796875, 54.56591796875, 
    57.56591796875, 60.56591796875, 63.56591796875, 66.56591796875, 
    69.56591796875, 72.56591796875, 75.56591796875, 78.56591796875, 
    81.56591796875, 84.56591796875, 87.56591796875, 90.56591796875,
  33.56591796875, 36.56591796875, 39.56591796875, 42.56591796875, 
    45.56591796875, 48.56591796875, 51.56591796875, 54.56591796875, 
    57.56591796875, 60.56591796875, 63.56591796875, 66.56591796875, 
    69.56591796875, 72.56591796875, 75.56591796875, 78.56591796875, 
    81.56591796875, 84.56591796875, 87.56591796875, 90.56591796875,
  30.29638671875, 33.29638671875, 36.29638671875, 39.29638671875, 
    42.29638671875, 45.29638671875, 48.29638671875, 51.29638671875, 
    54.29638671875, 57.29638671875, 60.29638671875, 63.29638671875, 
    66.29638671875, 69.29638671875, 72.29638671875, 75.29638671875, 
    78.29638671875, 81.29638671875, 84.29638671875, 87.29638671875,
  27.2783660888672, 30.2783660888672, 33.2783660888672, 36.2783660888672, 
    39.2783660888672, 42.2783660888672, 45.2783660888672, 48.2783660888672, 
    51.2783660888672, 54.2783660888672, 57.2783660888672, 60.2783660888672, 
    63.2783660888672, 66.2783660888672, 69.2783660888672, 72.2783660888672, 
    75.2783660888672, 78.2783660888672, 81.2783660888672, 84.2783660888672,
  24.2044448852539, 27.2044448852539, 30.2044448852539, 33.2044448852539, 
    36.2044448852539, 39.2044448852539, 42.2044448852539, 45.2044448852539, 
    48.2044448852539, 51.2044448852539, 54.2044448852539, 57.2044448852539, 
    60.2044448852539, 63.2044448852539, 66.2044448852539, 69.2044448852539, 
    72.2044448852539, 75.2044448852539, 78.2044448852539, 81.2044448852539,
  21.3540878295898, 24.3540878295898, 27.3540878295898, 30.3540878295898, 
    33.3540878295898, 36.3540878295898, 39.3540878295898, 42.3540878295898, 
    45.3540878295898, 48.3540878295898, 51.3540878295898, 54.3540878295898, 
    57.3540878295898, 60.3540878295898, 63.3540878295898, 66.3540878295898, 
    69.3540878295898, 72.3540878295898, 75.3540878295898, 78.3540878295898,
  18.2242889404297, 21.2242889404297, 24.2242889404297, 27.2242889404297, 
    30.2242889404297, 33.2242889404297, 36.2242889404297, 39.2242889404297, 
    42.2242889404297, 45.2242889404297, 48.2242889404297, 51.2242889404297, 
    54.2242889404297, 57.2242889404297, 60.2242889404297, 63.2242889404297, 
    66.2242889404297, 69.2242889404297, 72.2242889404297, 75.2242889404297,
  15.122428894043, 18.122428894043, 21.122428894043, 24.122428894043, 
    27.122428894043, 30.122428894043, 33.122428894043, 36.122428894043, 
    39.122428894043, 42.122428894043, 45.122428894043, 48.122428894043, 
    51.122428894043, 54.122428894043, 57.122428894043, 60.122428894043, 
    63.122428894043, 66.122428894043, 69.122428894043, 72.122428894043,
  11.824951171875, 14.824951171875, 17.824951171875, 20.824951171875, 
    23.824951171875, 26.824951171875, 29.824951171875, 32.824951171875, 
    35.824951171875, 38.824951171875, 41.824951171875, 44.824951171875, 
    47.824951171875, 50.824951171875, 53.824951171875, 56.824951171875, 
    59.824951171875, 62.824951171875, 65.824951171875, 68.824951171875,
  8.55542755126953, 11.5554275512695, 14.5554275512695, 17.5554275512695, 
    20.5554275512695, 23.5554275512695, 26.5554275512695, 29.5554275512695, 
    32.5554275512695, 35.5554275512695, 38.5554275512695, 41.5554275512695, 
    44.5554275512695, 47.5554275512695, 50.5554275512695, 53.5554275512695, 
    56.5554275512695, 59.5554275512695, 62.5554275512695, 65.5554275512695,
  8.55542755126953, 11.5554275512695, 14.5554275512695, 17.5554275512695, 
    20.5554275512695, 23.5554275512695, 26.5554275512695, 29.5554275512695, 
    32.5554275512695, 35.5554275512695, 38.5554275512695, 41.5554275512695, 
    44.5554275512695, 47.5554275512695, 50.5554275512695, 53.5554275512695, 
    56.5554275512695, 59.5554275512695, 62.5554275512695, 65.5554275512695,
  5.53739929199219, 8.53739929199219, 11.5373992919922, 14.5373992919922, 
    17.5373992919922, 20.5373992919922, 23.5373992919922, 26.5373992919922, 
    29.5373992919922, 32.5373992919922, 35.5373992919922, 38.5373992919922, 
    41.5373992919922, 44.5373992919922, 47.5373992919922, 50.5373992919922, 
    53.5373992919922, 56.5373992919922, 59.5373992919922, 62.5373992919922,
  2.26787185668945, 5.26787185668945, 8.26787185668945, 11.2678718566895, 
    14.2678718566895, 17.2678718566895, 20.2678718566895, 23.2678718566895, 
    26.2678718566895, 29.2678718566895, 32.2678718566895, 35.2678718566895, 
    38.2678718566895, 41.2678718566895, 44.2678718566895, 47.2678718566895, 
    50.2678718566895, 53.2678718566895, 56.2678718566895, 59.2678718566895,
  2.27779388427734, 5.27779388427734, 8.27779388427734, 11.2777938842773, 
    14.2777938842773, 17.2777938842773, 20.2777938842773, 23.2777938842773, 
    26.2777938842773, 29.2777938842773, 32.2777938842773, 35.2777938842773, 
    38.2777938842773, 41.2777938842773, 44.2777938842773, 47.2777938842773, 
    50.2777938842773, 53.2777938842773, 56.2777938842773, _,
  2.20387649536133, 5.20387649536133, 8.20387649536133, 11.2038764953613, 
    14.2038764953613, 17.2038764953613, 20.2038764953613, 23.2038764953613, 
    26.2038764953613, 29.2038764953613, 32.2038764953613, 35.2038764953613, 
    38.2038764953613, 41.2038764953613, 44.2038764953613, 47.2038764953613, 
    50.2038764953613, 53.2038764953613, _, _,
  1.96229553222656, 4.96229553222656, 7.96229553222656, 10.9622955322266, 
    13.9622955322266, 16.9622955322266, 19.9622955322266, 22.9622955322266, 
    25.9622955322266, 28.9622955322266, 31.9622955322266, 34.9622955322266, 
    37.9622955322266, 40.9622955322266, 43.9622955322266, 46.9622955322266, 
    49.9622955322266, _, _, _,
  1.88837814331055, 4.88837814331055, 7.88837814331055, 10.8883781433105, 
    13.8883781433105, 16.8883781433105, 19.8883781433105, 22.8883781433105, 
    25.8883781433105, 28.8883781433105, 31.8883781433105, 34.8883781433105, 
    37.8883781433105, 40.8883781433105, 43.8883781433105, 46.8883781433105, 
    _, _, _, _,
  1.73062896728516, 4.73062896728516, 7.73062896728516, 10.7306289672852, 
    13.7306289672852, 16.7306289672852, 19.7306289672852, 22.7306289672852, 
    25.7306289672852, 28.7306289672852, 31.7306289672852, 34.7306289672852, 
    37.7306289672852, 40.7306289672852, 43.7306289672852, _, _, _, _, _,
  1.79644012451172, 4.79644012451172, 7.79644012451172, 10.7964401245117, 
    13.7964401245117, 16.7964401245117, 19.7964401245117, 22.7964401245117, 
    25.7964401245117, 28.7964401245117, 31.7964401245117, 34.7964401245117, 
    37.7964401245117, 40.7964401245117, _, _, _, _, _, _,
  1.79644012451172, 4.79644012451172, 7.79644012451172, 10.7964401245117, 
    13.7964401245117, 16.7964401245117, 19.7964401245117, 22.7964401245117, 
    25.7964401245117, 28.7964401245117, 31.7964401245117, 34.7964401245117, 
    37.7964401245117, 40.7964401245117, _, _, _, _, _, _,
  1.55485534667969, 4.55485534667969, 7.55485534667969, 10.5548553466797, 
    13.5548553466797, 16.5548553466797, 19.5548553466797, 22.5548553466797, 
    25.5548553466797, 28.5548553466797, 31.5548553466797, 34.5548553466797, 
    37.5548553466797, _, _, _, _, _, _, _,
  1.62066650390625, 4.62066650390625, 7.62066650390625, 10.6206665039062, 
    13.6206665039062, 16.6206665039062, 19.6206665039062, 22.6206665039062, 
    25.6206665039062, 28.6206665039062, 31.6206665039062, 34.6206665039062, 
    _, _, _, _, _, _, _, _,
  1.40702629089355, 4.40702629089355, 7.40702629089355, 10.4070262908936, 
    13.4070262908936, 16.4070262908936, 19.4070262908936, 22.4070262908936, 
    25.4070262908936, 28.4070262908936, 31.4070262908936, _, _, _, _, _, _, 
    _, _, _,
  1.50078010559082, 4.50078010559082, 7.50078010559082, 10.5007801055908, 
    13.5007801055908, 16.5007801055908, 19.5007801055908, 22.5007801055908, 
    25.5007801055908, 28.5007801055908, _, _, _, _, _, _, _, _, _, _,
  1.45480918884277, 4.45480918884277, 7.45480918884277, 10.4548091888428, 
    13.4548091888428, 16.4548091888428, 19.4548091888428, 22.4548091888428, 
    25.4548091888428, _, _, _, _, _, _, _, _, _, _, _,
  1.5206184387207, 4.5206184387207, 7.5206184387207, 10.5206184387207, 
    13.5206184387207, 16.5206184387207, 19.5206184387207, 22.5206184387207, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  1.6423168182373, 4.6423168182373, 7.6423168182373, 10.6423168182373, 
    13.6423168182373, 16.6423168182373, 19.6423168182373, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  1.62429046630859, 4.62429046630859, 7.62429046630859, 10.6242904663086, 
    13.6242904663086, 16.6242904663086, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.62429046630859, 4.62429046630859, 7.62429046630859, 10.6242904663086, 
    13.6242904663086, 16.6242904663086, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.52243137359619, 4.52243137359619, 7.52243137359619, 10.5224313735962, 
    13.5224313735962, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.67207336425781, 4.67207336425781, 7.67207336425781, 10.6720733642578, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 echogram_sv =
  -31, -31, -31, -31, -31, -31, -31, -31, -31, -31, -31, -31, -31, -31, -31, 
    -31, -31, -31, -31, -31,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -67, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -67, -67, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -67, -61, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -61, -67, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -61, -67, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -55, -61, -61, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -67, -61, -61, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -61, -67, -61,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -61, -67, -61,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -67, -61,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -67, -73, -67,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -61,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, -73,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, -73, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, -73, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, -73, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    -73, _, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, 
    _, _, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, _, _, 
    _, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, _, _, 
    _, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, _, _, _, 
    _, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, _, _, _, _, _, 
    _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, _, _, _, _, _, _, _, 
    _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, -73, _, _, _, _, _, _, _, _, 
    _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, -73, _, _, _, _, _, _, _, _, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, -73, _, _, _, _, _, _, _, _, _, _, _, _,
  -73, -73, -73, -73, -73, -73, -73, _, _, _, _, _, _, _, _, _, _, _, _, _,
  -73, -73, -73, -73, -73, -73, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  -73, -73, -73, -73, -73, -73, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  -73, -55, -61, -73, -73, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  -67, -31, -73, -73, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 lat = 59.8421046403177, 59.8419970771558, 59.8419375741301, 
    59.8418986683056, 59.8418506081694, 59.8418071251891, 59.8417636422088, 
    59.8417224478064, 59.8416766762481, 59.8416354818457, 59.8415919988654, 
    59.8415508044629, 59.8415050329047, 59.8414615499244, 59.841418066944, 
    59.8413768725416, 59.8413311009834, 59.841287618003, 59.8412487121785, 
    59.8412029406203, 59.8411594576399, 59.8411159746596, 59.8410747802572, 
    59.8410312972768, 59.8409878142965, 59.8409420427383, 59.8409008483359, 
    59.8408596539334, 59.8408138823752, 59.8407703993949, 59.8407292049924, 
    59.8406857220121, 59.8406422390318, 59.8405964674735, 59.8405552730711, 
    59.8405117900908, 59.8404683071104, 59.8404248241301, 59.8403813411498, 
    59.8403401467474, 59.8402989523449, 59.8402508922088, 59.8402096978064, 
    59.840166214826, 59.8401227318457, 59.8400792488654, 59.840035765885, 
    59.8399922829047, 59.8399510885023, 59.8399098940998, 59.8398618339637, 
    59.8398206395613, 59.8397771565809, 59.8397359621785, 59.8396901906203, 
    59.8396467076399, 59.8396055132375, 59.8395620302572, 59.8395208358548, 
    59.8394750642965, 59.8394315813162, 59.8393880983359, 59.8393469039334, 
    59.8393011323752, 59.8392576493949, 59.8392164549924 ;

 lon = -149.475288063162, -149.475348910741, -149.475382571104, 
    -149.475404579803, -149.47543176702, -149.475456364977, 
    -149.475480962935, -149.475504266263, -149.47553015885, 
    -149.475553462179, -149.475578060136, -149.475601363464, 
    -149.475627256051, -149.475651854009, -149.475676451967, 
    -149.475699755295, -149.475725647882, -149.47575024584, 
    -149.475772254539, -149.475798147126, -149.475822745083, 
    -149.475847343041, -149.475870646369, -149.475895244327, 
    -149.475919842284, -149.475945734871, -149.4759690382, -149.475992341528, 
    -149.476018234115, -149.476042832073, -149.476066135401, 
    -149.476090733359, -149.476115331316, -149.476141223903, 
    -149.476164527231, -149.476189125189, -149.476213723147, 
    -149.476238321104, -149.476262919062, -149.47628622239, 
    -149.476309525719, -149.476336712935, -149.476360016263, 
    -149.476384614221, -149.476409212179, -149.476433810136, 
    -149.476458408094, -149.476483006051, -149.47650630938, 
    -149.476529612708, -149.476556799924, -149.476580103253, 
    -149.47660470121, -149.476628004539, -149.476653897126, 
    -149.476678495083, -149.476701798411, -149.476726396369, 
    -149.476749699697, -149.476775592284, -149.476800190242, -149.4768247882, 
    -149.476848091528, -149.476873984115, -149.476898582073, -149.476921885401 ;

 lat_uv = _ ;

 lon_uv = _ ;

 time_uv = _ ;

 profile_id = 1710362769 ;

 profile_lat = 59.840776394132 ;

 profile_lon = -149.4760394409 ;

 profile_time = 1079211350.06525 ;

 u = _ ;

 v = _ ;

 platform = _ ;

 instrument_ctd = _ ;

 trajectory = "unit_507-20240304T0000" ;
}
